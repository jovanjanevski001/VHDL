library ieee;
use ieee.std_logic_1164.all;

package decoder7seg_package is 
	
	constant	c_0	:	std_logic_vector(6 downto 0)	:= "1000000";
	constant	c_1	:	std_logic_vector(6 downto 0)	:= "1111001";
	constant	c_2	:	std_logic_vector(6 downto 0)	:= "0100100";
	constant	c_3	:	std_logic_vector(6 downto 0)	:= "0110000";
	constant	c_4	:	std_logic_vector(6 downto 0)	:= "0011001";
	constant	c_5	:	std_logic_vector(6 downto 0)	:= "0010010";
	constant	c_6	:	std_logic_vector(6 downto 0)	:= "0000010";
	constant	c_7	:	std_logic_vector(6 downto 0)	:= "1111000";
	constant	c_8	:	std_logic_vector(6 downto 0)	:= "0000000";
	constant	c_9	:	std_logic_vector(6 downto 0)	:= "0011000";
	constant	c_A	:	std_logic_vector(6 downto 0)	:= "0001000";
	constant	c_B	:	std_logic_vector(6 downto 0)	:= "0000011";
	constant	c_C	:	std_logic_vector(6 downto 0)	:= "0100111";
	constant	c_D	:	std_logic_vector(6 downto 0)	:= "0100001";
	constant	c_E	:	std_logic_vector(6 downto 0)	:= "0000110";
	constant	c_F	:	std_logic_vector(6 downto 0)	:= "0001110";
	
end package decoder7seg_package;

package body decoder7seg_package is
end package body decoder7seg_package;